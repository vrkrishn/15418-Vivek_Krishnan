module decision_tree
    #(parameter S, parameter dataSize)
    input logic 
